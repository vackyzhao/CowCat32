module tb_CPU();
SynCPU sim_CPU();
endmodule