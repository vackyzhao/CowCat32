
// font_rom.v
// 字符点阵ROM模块，用于存储字符0-9和a-z的8x8点阵数据
module font_rom(
    input wire [7:0] ascii_code,  // ASCII码输入
    input wire [2:0] row,         // 行号输入 (0-7)
    output reg [7:0] data         // 输出当前行的点阵数据
);
// 字符 0-9 的 8x8 点阵
reg [7:0] font [48:122][0:7]; // ASCII 码 48-57 对应 0-9

initial begin
    // Character '0' ASCII 48
font[8'h30][0] = 8'b00000000;
font[8'h30][1] = 8'b00000000;
font[8'h30][2] = 8'b01110000;
font[8'h30][3] = 8'b11011000;
font[8'h30][4] = 8'b11011000;
font[8'h30][5] = 8'b11011000;
font[8'h30][6] = 8'b11011000;
font[8'h30][7] = 8'b11011000;

// Character '1' ASCII 49
font[8'h31][0] = 8'b00000000;
font[8'h31][1] = 8'b00000000;
font[8'h31][2] = 8'b00110000;
font[8'h31][3] = 8'b11110000;
font[8'h31][4] = 8'b00110000;
font[8'h31][5] = 8'b00110000;
font[8'h31][6] = 8'b00110000;
font[8'h31][7] = 8'b00110000;

// Character '2' ASCII 50
font[8'h32][0] = 8'b00000000;
font[8'h32][1] = 8'b00000000;
font[8'h32][2] = 8'b01110000;
font[8'h32][3] = 8'b11011000;
font[8'h32][4] = 8'b00011000;
font[8'h32][5] = 8'b00110000;
font[8'h32][6] = 8'b01100000;
font[8'h32][7] = 8'b11011000;

// Character '3' ASCII 51
font[8'h33][0] = 8'b00000000;
font[8'h33][1] = 8'b00000000;
font[8'h33][2] = 8'b01110000;
font[8'h33][3] = 8'b11011000;
font[8'h33][4] = 8'b00011000;
font[8'h33][5] = 8'b01110000;
font[8'h33][6] = 8'b00011000;
font[8'h33][7] = 8'b11011000;

// Character '4' ASCII 52
font[8'h34][0] = 8'b00000000;
font[8'h34][1] = 8'b00000000;
font[8'h34][2] = 8'b00011000;
font[8'h34][3] = 8'b00111000;
font[8'h34][4] = 8'b01011000;
font[8'h34][5] = 8'b11011000;
font[8'h34][6] = 8'b11111100;
font[8'h34][7] = 8'b00011000;

// Character '5' ASCII 53
font[8'h35][0] = 8'b00000000;
font[8'h35][1] = 8'b00000000;
font[8'h35][2] = 8'b11111000;
font[8'h35][3] = 8'b11000000;
font[8'h35][4] = 8'b11110000;
font[8'h35][5] = 8'b11011000;
font[8'h35][6] = 8'b00011000;
font[8'h35][7] = 8'b10011000;

// Character '6' ASCII 54
font[8'h36][0] = 8'b00000000;
font[8'h36][1] = 8'b00000000;
font[8'h36][2] = 8'b01110000;
font[8'h36][3] = 8'b11011000;
font[8'h36][4] = 8'b11000000;
font[8'h36][5] = 8'b11110000;
font[8'h36][6] = 8'b11011000;
font[8'h36][7] = 8'b11011000;

// Character '7' ASCII 55
font[8'h37][0] = 8'b00000000;
font[8'h37][1] = 8'b00000000;
font[8'h37][2] = 8'b11111000;
font[8'h37][3] = 8'b11011000;
font[8'h37][4] = 8'b00011000;
font[8'h37][5] = 8'b00110000;
font[8'h37][6] = 8'b00110000;
font[8'h37][7] = 8'b01100000;

// Character '8' ASCII 56
font[8'h38][0] = 8'b00000000;
font[8'h38][1] = 8'b00000000;
font[8'h38][2] = 8'b01110000;
font[8'h38][3] = 8'b11011000;
font[8'h38][4] = 8'b11011000;
font[8'h38][5] = 8'b01110000;
font[8'h38][6] = 8'b11011000;
font[8'h38][7] = 8'b11011000;

// Character '9' ASCII 57
font[8'h39][0] = 8'b00000000;
font[8'h39][1] = 8'b00000000;
font[8'h39][2] = 8'b01110000;
font[8'h39][3] = 8'b11011000;
font[8'h39][4] = 8'b11011000;
font[8'h39][5] = 8'b01111000;
font[8'h39][6] = 8'b00011000;
font[8'h39][7] = 8'b11011000;

// Character 'a' ASCII 97
font[8'h61][0] = 8'b00000000;
font[8'h61][1] = 8'b00000000;
font[8'h61][2] = 8'b00000000;
font[8'h61][3] = 8'b00000000;
font[8'h61][4] = 8'b01110000;
font[8'h61][5] = 8'b11011000;
font[8'h61][6] = 8'b01111000;
font[8'h61][7] = 8'b11011000;

// Character 'b' ASCII 98
font[8'h62][0] = 8'b00000000;
font[8'h62][1] = 8'b00000000;
font[8'h62][2] = 8'b11000000;
font[8'h62][3] = 8'b11000000;
font[8'h62][4] = 8'b11110000;
font[8'h62][5] = 8'b11011000;
font[8'h62][6] = 8'b11011000;
font[8'h62][7] = 8'b11011000;

// Character 'c' ASCII 99
font[8'h63][0] = 8'b00000000;
font[8'h63][1] = 8'b00000000;
font[8'h63][2] = 8'b00000000;
font[8'h63][3] = 8'b00000000;
font[8'h63][4] = 8'b01110000;
font[8'h63][5] = 8'b11011000;
font[8'h63][6] = 8'b11000000;
font[8'h63][7] = 8'b11011000;

// Character 'd' ASCII 100
font[8'h64][0] = 8'b00000000;
font[8'h64][1] = 8'b00000000;
font[8'h64][2] = 8'b00111000;
font[8'h64][3] = 8'b00011000;
font[8'h64][4] = 8'b01111000;
font[8'h64][5] = 8'b11011000;
font[8'h64][6] = 8'b11011000;
font[8'h64][7] = 8'b11011000;

// Character 'e' ASCII 101
font[8'h65][0] = 8'b00000000;
font[8'h65][1] = 8'b00000000;
font[8'h65][2] = 8'b00000000;
font[8'h65][3] = 8'b00000000;
font[8'h65][4] = 8'b01110000;
font[8'h65][5] = 8'b11011000;
font[8'h65][6] = 8'b11111000;
font[8'h65][7] = 8'b11000000;

// Character 'f' ASCII 102
font[8'h66][0] = 8'b00000000;
font[8'h66][1] = 8'b00000000;
font[8'h66][2] = 8'b00111000;
font[8'h66][3] = 8'b01100000;
font[8'h66][4] = 8'b11111000;
font[8'h66][5] = 8'b01100000;
font[8'h66][6] = 8'b01100000;
font[8'h66][7] = 8'b01100000;

// Character 'g' ASCII 103
font[8'h67][0] = 8'b00000000;
font[8'h67][1] = 8'b00000000;
font[8'h67][2] = 8'b00000000;
font[8'h67][3] = 8'b00000000;
font[8'h67][4] = 8'b01101100;
font[8'h67][5] = 8'b11011000;
font[8'h67][6] = 8'b11011000;
font[8'h67][7] = 8'b11011000;

// Character 'h' ASCII 104
font[8'h68][0] = 8'b00000000;
font[8'h68][1] = 8'b00000000;
font[8'h68][2] = 8'b11000000;
font[8'h68][3] = 8'b11000000;
font[8'h68][4] = 8'b11110000;
font[8'h68][5] = 8'b11011000;
font[8'h68][6] = 8'b11011000;
font[8'h68][7] = 8'b11011000;

// Character 'i' ASCII 105
font[8'h69][0] = 8'b00000000;
font[8'h69][1] = 8'b00000000;
font[8'h69][2] = 8'b00110000;
font[8'h69][3] = 8'b00000000;
font[8'h69][4] = 8'b11110000;
font[8'h69][5] = 8'b00110000;
font[8'h69][6] = 8'b00110000;
font[8'h69][7] = 8'b00110000;

// Character 'j' ASCII 106
font[8'h6A][0] = 8'b00000000;
font[8'h6A][1] = 8'b00000000;
font[8'h6A][2] = 8'b00110000;
font[8'h6A][3] = 8'b00000000;
font[8'h6A][4] = 8'b11110000;
font[8'h6A][5] = 8'b00110000;
font[8'h6A][6] = 8'b00110000;
font[8'h6A][7] = 8'b00110000;

// Character 'k' ASCII 107
font[8'h6B][0] = 8'b00000000;
font[8'h6B][1] = 8'b00000000;
font[8'h6B][2] = 8'b11000000;
font[8'h6B][3] = 8'b11000000;
font[8'h6B][4] = 8'b11011000;
font[8'h6B][5] = 8'b11110000;
font[8'h6B][6] = 8'b11100000;
font[8'h6B][7] = 8'b11110000;

// Character 'l' ASCII 108
font[8'h6C][0] = 8'b00000000;
font[8'h6C][1] = 8'b00000000;
font[8'h6C][2] = 8'b11110000;
font[8'h6C][3] = 8'b00110000;
font[8'h6C][4] = 8'b00110000;
font[8'h6C][5] = 8'b00110000;
font[8'h6C][6] = 8'b00110000;
font[8'h6C][7] = 8'b00110000;

// Character 'm' ASCII 109
font[8'h6D][0] = 8'b00000000;
font[8'h6D][1] = 8'b00000000;
font[8'h6D][2] = 8'b00000000;
font[8'h6D][3] = 8'b00000000;
font[8'h6D][4] = 8'b11110000;
font[8'h6D][5] = 8'b11111000;
font[8'h6D][6] = 8'b10101000;
font[8'h6D][7] = 8'b10101000;

// Character 'n' ASCII 110
font[8'h6E][0] = 8'b00000000;
font[8'h6E][1] = 8'b00000000;
font[8'h6E][2] = 8'b00000000;
font[8'h6E][3] = 8'b00000000;
font[8'h6E][4] = 8'b10110000;
font[8'h6E][5] = 8'b11011000;
font[8'h6E][6] = 8'b11011000;
font[8'h6E][7] = 8'b11011000;

// Character 'o' ASCII 111
font[8'h6F][0] = 8'b00000000;
font[8'h6F][1] = 8'b00000000;
font[8'h6F][2] = 8'b00000000;
font[8'h6F][3] = 8'b00000000;
font[8'h6F][4] = 8'b01110000;
font[8'h6F][5] = 8'b11011000;
font[8'h6F][6] = 8'b11011000;
font[8'h6F][7] = 8'b11011000;

// Character 'p' ASCII 112
font[8'h70][0] = 8'b00000000;
font[8'h70][1] = 8'b00000000;
font[8'h70][2] = 8'b00000000;
font[8'h70][3] = 8'b00000000;
font[8'h70][4] = 8'b11110000;
font[8'h70][5] = 8'b11011000;
font[8'h70][6] = 8'b11011000;
font[8'h70][7] = 8'b11011000;

// Character 'q' ASCII 113
font[8'h71][0] = 8'b00000000;
font[8'h71][1] = 8'b00000000;
font[8'h71][2] = 8'b00000000;
font[8'h71][3] = 8'b00000000;
font[8'h71][4] = 8'b01101100;
font[8'h71][5] = 8'b11011000;
font[8'h71][6] = 8'b11011000;
font[8'h71][7] = 8'b11011000;

// Character 'r' ASCII 114
font[8'h72][0] = 8'b00000000;
font[8'h72][1] = 8'b00000000;
font[8'h72][2] = 8'b00000000;
font[8'h72][3] = 8'b00000000;
font[8'h72][4] = 8'b11011100;
font[8'h72][5] = 8'b01110100;
font[8'h72][6] = 8'b01100000;
font[8'h72][7] = 8'b01100000;

// Character 's' ASCII 115
font[8'h73][0] = 8'b00000000;
font[8'h73][1] = 8'b00000000;
font[8'h73][2] = 8'b00000000;
font[8'h73][3] = 8'b00000000;
font[8'h73][4] = 8'b01111000;
font[8'h73][5] = 8'b11100000;
font[8'h73][6] = 8'b01111000;
font[8'h73][7] = 8'b00011100;

// Character 't' ASCII 116
font[8'h74][0] = 8'b00000000;
font[8'h74][1] = 8'b00000000;
font[8'h74][2] = 8'b01100000;
font[8'h74][3] = 8'b01100000;
font[8'h74][4] = 8'b11111000;
font[8'h74][5] = 8'b01100000;
font[8'h74][6] = 8'b01100000;
font[8'h74][7] = 8'b01101100;

// Character 'u' ASCII 117
font[8'h75][0] = 8'b00000000;
font[8'h75][1] = 8'b00000000;
font[8'h75][2] = 8'b00000000;
font[8'h75][3] = 8'b00000000;
font[8'h75][4] = 8'b11011000;
font[8'h75][5] = 8'b11011000;
font[8'h75][6] = 8'b11011000;
font[8'h75][7] = 8'b11011000;

// Character 'v' ASCII 118
font[8'h76][0] = 8'b00000000;
font[8'h76][1] = 8'b00000000;
font[8'h76][2] = 8'b00000000;
font[8'h76][3] = 8'b00000000;
font[8'h76][4] = 8'b11011000;
font[8'h76][5] = 8'b11011000;
font[8'h76][6] = 8'b01110000;
font[8'h76][7] = 8'b01110000;

// Character 'w' ASCII 119
font[8'h77][0] = 8'b00000000;
font[8'h77][1] = 8'b00000000;
font[8'h77][2] = 8'b00000000;
font[8'h77][3] = 8'b00000000;
font[8'h77][4] = 8'b10101100;
font[8'h77][5] = 8'b10101000;
font[8'h77][6] = 8'b11111000;
font[8'h77][7] = 8'b01111000;

// Character 'x' ASCII 120
font[8'h78][0] = 8'b00000000;
font[8'h78][1] = 8'b00000000;
font[8'h78][2] = 8'b00000000;
font[8'h78][3] = 8'b00000000;
font[8'h78][4] = 8'b11101100;
font[8'h78][5] = 8'b01111000;
font[8'h78][6] = 8'b00110000;
font[8'h78][7] = 8'b01111000;

// Character 'y' ASCII 121
font[8'h79][0] = 8'b00000000;
font[8'h79][1] = 8'b00000000;
font[8'h79][2] = 8'b00000000;
font[8'h79][3] = 8'b00000000;
font[8'h79][4] = 8'b11011100;
font[8'h79][5] = 8'b11011000;
font[8'h79][6] = 8'b11011000;
font[8'h79][7] = 8'b01010000;

// Character 'z' ASCII 122
font[8'h7A][0] = 8'b00000000;
font[8'h7A][1] = 8'b00000000;
font[8'h7A][2] = 8'b00000000;
font[8'h7A][3] = 8'b00000000;
font[8'h7A][4] = 8'b11111000;
font[8'h7A][5] = 8'b10110000;
font[8'h7A][6] = 8'b01100000;
font[8'h7A][7] = 8'b11011000;


end

   // 根据输入的ASCII码和行号输出对应的字符点阵行数据
    always @(*) begin
        if (ascii_code >= 8'h30 && ascii_code <= 8'h39 || ascii_code >= 8'h61 && ascii_code <= 8'h7A) begin
            data = font[ascii_code][row];
        end else begin
            data = 8'b00000000;  // 不在范围内时输出空白行
        end
    end

endmodule